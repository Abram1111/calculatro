//Top Level Entity
module Calculator(SW,HEX00,HEX01,HEX02,HEX03,HEX04,HEX05,HEX06,HEX10,HEX11,HEX12,HEX13,HEX14,HEX15,HEX16);
	input [7:0] SW;
	output HEX00,HEX01,HEX02,HEX03,HEX04,HEX05,HEX06,HEX10,HEX11,HEX12,HEX13,HEX14,HEX15,HEX16;
	
	wire [4:0] sum;
	
	four_ripple_adder mainadder(SW[3:0],SW[7:4],sum);
	segment_display maindisplay(sum,HEX00,HEX01,HEX02,HEX03,HEX04,HEX05,HEX06,HEX10,HEX11,HEX12,HEX13,HEX14,HEX15,HEX16);

endmodule
